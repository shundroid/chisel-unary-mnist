`define WIDTH 3
module baseline(input clock, output io_out);
logic [WIDTH-1:0] mul1;

endmodule